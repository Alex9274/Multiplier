--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   00:35:30 01/09/2015
-- Design Name:   
-- Module Name:   C:/Users/Alex/Desktop/2.5.1/Top_tb.vhd
-- Project Name:  Multiplicador_8_bits
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: TOP
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Top_tb IS
END Top_tb;
 
ARCHITECTURE behavior OF Top_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT TOP
    PORT(
         reset : IN  std_logic;
         clk : IN  std_logic;
         din : IN  std_logic_vector(7 downto 0);
         enter : IN  std_logic;
         segments : OUT  std_logic_vector(6 downto 0);
         digits : OUT  std_logic_vector(3 downto 0);
         signo : OUT  std_logic;
         overflow : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal reset : std_logic;-- := '0';
   signal clk : std_logic;-- := '0';
   signal din : std_logic_vector(7 downto 0);-- := (others => '0');
   signal enter : std_logic := '0';

 	--Outputs
   signal segments : std_logic_vector(6 downto 0);
   signal digits : std_logic_vector(3 downto 0);
   signal signo : std_logic;
   signal overflow : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: TOP PORT MAP (
          reset => reset,
          clk => clk,
          din => din,
          enter => enter,
          segments => segments,
          digits => digits,
          signo => signo,
          overflow => overflow
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 50 ns;	

      --wait for clk_period*10;

      -- insert stimulus here 
		
		
		enter <= '1';			--Pulsamos enter 	
		--wait for 1 ns;
		enter <= '0';
		din <= "00000010";	--Metemos primer n�mero
		
		
		enter <= '1';			--Pulsamos enter
		wait for 50 ns;
		enter <= '0';
		din <= "10111101";	--Metemos segundo n�mero
		
		wait for 20 ns;
		enter <= '1';			--Pulsamos enter para multiplicar
		wait for 5 ns;
		enter <= '0';
		
		wait for 50 ns;
		
		
		
		
     
   end process;

END;
