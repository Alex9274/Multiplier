`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:16:48 01/04/2015 
// Design Name: 
// Module Name:    Conv_14 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Conv_14(
    input din14,
    output dout1,
    output dout2,
    output dout3,
    output dout4,
    output dout
    );


endmodule
